* TLE2082 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 04/06/94 AT 15:13
* REV N/A        SUPPLIES +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLE2082  1 2 3 4 5
*
  C1   11 12 1.2E-12
  C2    6  7 10.00E-12
  CPSR 85 86 159E-9
  DCM+ 81 82 DX
  DCM- 83 81 DX
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  ECMR 84 99 (2,99) 1
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  EPSR 85 0 POLY(1) (3,4) -336E-6 11.2E-6
  ENSE 89 2 POLY(1) (88,0) 490E-6 1
  FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 5.607E6 -6E6 6E6 6E6 -6E6 37.8E6
  GA    6  0 11 12 333.0E-6
  GCM 0  6 10 99 7.436E-9
  GPSR 85 86 (85,86) 100E-6
  GRD1 60 11 (60,11) 333E-6
  GRD2 60 12 (60,12) 333E-6
  HLIM 90  0 VLIM 1K
  HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
  IRP 3 4 1.3E-3
  ISS   3 10 DC 400.0E-6
  IIO 2 0 6E-12
  I1 88 0 1E-21
  J1   11  89 10 JX
  J2   12  80 10 JX
  R2    6  9 100.0E3
  RCM 84 81 1K
  RN1 88 0 8000
  RO1   8  5 80
  RO2   7 99 80
  RSS  10 99 500.0E3
  VAD 60 4 -.6
  VCM+ 82 99 14.4
  VCM- 83 99 -11.3
  VB    9  0 DC 0
  VC 3 53 DC 1.7
  VE   54  4 DC 1.7
  VLIM  7  8 DC 0
  VLP  91  0 DC 45
  VLN   0 92 DC 45
  VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=554.5E-6 VTO=-.564 KF=7E-18)
.ENDS

